assign strg_ub_agg_read_addr_gen_0_starting_addr = 0;
assign strg_ub_input_addr_gen_starting_addr = 0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr = 4;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality = 3;
assign strg_ub_loops_in2buf_autovec_write_dimensionality = 3;
assign strg_ub_output_addr_gen_starting_addr = 0;
assign strg_ub_tb_write_addr_gen_0_starting_addr = 0;
assign strg_ub_tb_write_addr_gen_1_starting_addr = 0;
assign strg_ub_out_port_sel_addr_starting_addr = 0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr = 29;
assign loops_buf2out_autovec_read_dimensionality = 4;
assign strg_ub_loops_buf2out_out_sel_dimensionality = 4;
assign strg_ub_agg_write_addr_gen_0_starting_addr = 0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr = 0;
assign strg_ub_loops_in2buf_0_dimensionality = 3;
assign strg_ub_tb_read_addr_gen_0_starting_addr = 0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr = 32;
assign strg_ub_loops_buf2out_read_0_dimensionality = 3;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality = 3;
assign strg_ub_tb_read_addr_gen_1_starting_addr = 16;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr = 32;
assign strg_ub_loops_buf2out_read_1_dimensionality = 3;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality = 3;
assign chain_idx_input = 0;
assign chain_idx_output = 0;
assign enable_chain_input = 0;
assign enable_chain_output = 0;
assign chain_valid_in_reg_sel = 1;
assign chain_valid_in_reg_value = 0;
assign flush_reg_sel = 1;
assign flush_reg_value = 0;
assign ren_in_reg_sel = 1;
assign ren_in_reg_value = 0;
assign wen_in_reg_sel = 1;
assign wen_in_reg_value = 0;
assign mode = 0;
assign tile_en = 1;
assign strg_ub_loops_in2buf_0_ranges[0] = 2;
assign strg_ub_agg_write_addr_gen_0_strides[0] = 1;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[0] = 1;
assign strg_ub_loops_in2buf_0_ranges[1] = 30;
assign strg_ub_agg_write_addr_gen_0_strides[1] = -3;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[1] = 1;
assign strg_ub_loops_in2buf_0_ranges[2] = -1;
assign strg_ub_agg_write_addr_gen_0_strides[2] = -3;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[2] = -127;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[0] = 2;
assign strg_ub_agg_read_addr_gen_0_strides[0] = 4;
assign strg_ub_loops_in2buf_autovec_write_ranges[0] = 2;
assign strg_ub_input_addr_gen_strides[0] = 1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[0] = 4;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[1] = 6;
assign strg_ub_agg_read_addr_gen_0_strides[1] = 4;
assign strg_ub_loops_in2buf_autovec_write_ranges[1] = 6;
assign strg_ub_input_addr_gen_strides[1] = 1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[1] = 4;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[2] = -1;
assign strg_ub_agg_read_addr_gen_0_strides[2] = -124;
assign strg_ub_loops_in2buf_autovec_write_ranges[2] = -1;
assign strg_ub_input_addr_gen_strides[2] = -31;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[2] = -124;
assign strg_ub_loops_buf2out_autovec_read_ranges[0] = 0;
assign strg_ub_output_addr_gen_strides[0] = 4;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[0] = 2;
assign strg_ub_loops_buf2out_out_sel_ranges[0] = 0;
assign strg_ub_out_port_sel_addr_strides[0] = 1;
assign strg_ub_tb_write_addr_gen_0_strides[0] = 1;
assign strg_ub_tb_write_addr_gen_1_strides[0] = 1;
assign strg_ub_loops_buf2out_autovec_read_ranges[1] = 2;
assign strg_ub_output_addr_gen_strides[1] = -3;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[1] = 2;
assign strg_ub_loops_buf2out_out_sel_ranges[1] = 2;
assign strg_ub_out_port_sel_addr_strides[1] = -1;
assign strg_ub_tb_write_addr_gen_0_strides[1] = -1;
assign strg_ub_tb_write_addr_gen_1_strides[1] = -1;
assign strg_ub_loops_buf2out_autovec_read_ranges[2] = 4;
assign strg_ub_output_addr_gen_strides[2] = -3;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[2] = 2;
assign strg_ub_loops_buf2out_out_sel_ranges[2] = 4;
assign strg_ub_out_port_sel_addr_strides[2] = -1;
assign strg_ub_tb_write_addr_gen_0_strides[2] = -1;
assign strg_ub_tb_write_addr_gen_1_strides[2] = -1;
assign strg_ub_loops_buf2out_autovec_read_ranges[3] = -1;
assign strg_ub_output_addr_gen_strides[3] = -27;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[3] = -94;
assign strg_ub_loops_buf2out_out_sel_ranges[3] = -1;
assign strg_ub_out_port_sel_addr_strides[3] = -1;
assign strg_ub_tb_write_addr_gen_0_strides[3] = -1;
assign strg_ub_tb_write_addr_gen_1_strides[3] = -1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[0] = 14;
assign strg_ub_loops_buf2out_read_0_ranges[0] = 14;
assign strg_ub_tb_read_addr_gen_0_strides[0] = 1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[0] = 1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[1] = 4;
assign strg_ub_loops_buf2out_read_0_ranges[1] = 4;
assign strg_ub_tb_read_addr_gen_0_strides[1] = 1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[1] = 1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[2] = -1;
assign strg_ub_loops_buf2out_read_0_ranges[2] = -1;
assign strg_ub_tb_read_addr_gen_0_strides[2] = -95;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[2] = -95;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[0] = 14;
assign strg_ub_loops_buf2out_read_1_ranges[0] = 14;
assign strg_ub_tb_read_addr_gen_1_strides[0] = 1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[0] = 1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[1] = 4;
assign strg_ub_loops_buf2out_read_1_ranges[1] = 4;
assign strg_ub_tb_read_addr_gen_1_strides[1] = 1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[1] = 1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[2] = -1;
assign strg_ub_loops_buf2out_read_1_ranges[2] = -1;
assign strg_ub_tb_read_addr_gen_1_strides[2] = -95;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[2] = -95;

assign strg_ub_agg_read_addr_gen_0_starting_addr = 'd0;
assign strg_ub_input_addr_gen_starting_addr = 'd0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr = 'd4;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality = 'd3;
assign strg_ub_loops_in2buf_autovec_write_dimensionality = 'd3;
assign strg_ub_output_addr_gen_starting_addr = 'd0;
assign strg_ub_tb_write_addr_gen_0_starting_addr = 'd0;
assign strg_ub_tb_write_addr_gen_1_starting_addr = 'd0;
assign strg_ub_out_port_sel_addr_starting_addr = 'd0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr = 'd29;
assign loops_buf2out_autovec_read_dimensionality = 'd4;
assign strg_ub_loops_buf2out_out_sel_dimensionality = 'd4;
assign strg_ub_agg_write_addr_gen_0_starting_addr = 'd0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr = 'd0;
assign strg_ub_loops_in2buf_0_dimensionality = 'd3;
assign strg_ub_tb_read_addr_gen_0_starting_addr = 'd0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr = 'd32;
assign strg_ub_loops_buf2out_read_0_dimensionality = 'd3;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality = 'd3;
assign strg_ub_tb_read_addr_gen_1_starting_addr = 'd16;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr = 'd32;
assign strg_ub_loops_buf2out_read_1_dimensionality = 'd3;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality = 'd3;
assign chain_idx_input = 'd0;
assign chain_idx_output = 'd0;
assign enable_chain_input = 'd0;
assign enable_chain_output = 'd0;
assign chain_valid_in_reg_sel = 'd1;
assign chain_valid_in_reg_value = 'd0;
assign flush_reg_sel = 'd1;
assign flush_reg_value = 'd0;
assign ren_in_reg_sel = 'd1;
assign ren_in_reg_value = 'd0;
assign wen_in_reg_sel = 'd1;
assign wen_in_reg_value = 'd0;
assign mode = 'd0;
assign tile_en = 'd1;
assign strg_ub_loops_in2buf_0_ranges[0] = 'd2;
assign strg_ub_agg_write_addr_gen_0_strides[0] = 'd1;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[0] = 'd1;
assign strg_ub_loops_in2buf_0_ranges[1] = 'd30;
assign strg_ub_agg_write_addr_gen_0_strides[1] = 'd-3;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[1] = 'd1;
assign strg_ub_loops_in2buf_0_ranges[2] = 'd-1;
assign strg_ub_agg_write_addr_gen_0_strides[2] = 'd-3;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[2] = 'd-127;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[0] = 'd2;
assign strg_ub_agg_read_addr_gen_0_strides[0] = 'd4;
assign strg_ub_loops_in2buf_autovec_write_ranges[0] = 'd2;
assign strg_ub_input_addr_gen_strides[0] = 'd1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[0] = 'd4;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[1] = 'd6;
assign strg_ub_agg_read_addr_gen_0_strides[1] = 'd4;
assign strg_ub_loops_in2buf_autovec_write_ranges[1] = 'd6;
assign strg_ub_input_addr_gen_strides[1] = 'd1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[1] = 'd4;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[2] = 'd-1;
assign strg_ub_agg_read_addr_gen_0_strides[2] = 'd-124;
assign strg_ub_loops_in2buf_autovec_write_ranges[2] = 'd-1;
assign strg_ub_input_addr_gen_strides[2] = 'd-31;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[2] = 'd-124;
assign strg_ub_loops_buf2out_autovec_read_ranges[0] = 'd0;
assign strg_ub_output_addr_gen_strides[0] = 'd4;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[0] = 'd2;
assign strg_ub_loops_buf2out_out_sel_ranges[0] = 'd0;
assign strg_ub_out_port_sel_addr_strides[0] = 'd1;
assign strg_ub_tb_write_addr_gen_0_strides[0] = 'd1;
assign strg_ub_tb_write_addr_gen_1_strides[0] = 'd1;
assign strg_ub_loops_buf2out_autovec_read_ranges[1] = 'd2;
assign strg_ub_output_addr_gen_strides[1] = 'd-3;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[1] = 'd2;
assign strg_ub_loops_buf2out_out_sel_ranges[1] = 'd2;
assign strg_ub_out_port_sel_addr_strides[1] = 'd-1;
assign strg_ub_tb_write_addr_gen_0_strides[1] = 'd-1;
assign strg_ub_tb_write_addr_gen_1_strides[1] = 'd-1;
assign strg_ub_loops_buf2out_autovec_read_ranges[2] = 'd4;
assign strg_ub_output_addr_gen_strides[2] = 'd-3;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[2] = 'd2;
assign strg_ub_loops_buf2out_out_sel_ranges[2] = 'd4;
assign strg_ub_out_port_sel_addr_strides[2] = 'd-1;
assign strg_ub_tb_write_addr_gen_0_strides[2] = 'd-1;
assign strg_ub_tb_write_addr_gen_1_strides[2] = 'd-1;
assign strg_ub_loops_buf2out_autovec_read_ranges[3] = 'd-1;
assign strg_ub_output_addr_gen_strides[3] = 'd-27;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[3] = 'd-94;
assign strg_ub_loops_buf2out_out_sel_ranges[3] = 'd-1;
assign strg_ub_out_port_sel_addr_strides[3] = 'd-1;
assign strg_ub_tb_write_addr_gen_0_strides[3] = 'd-1;
assign strg_ub_tb_write_addr_gen_1_strides[3] = 'd-1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[0] = 'd14;
assign strg_ub_loops_buf2out_read_0_ranges[0] = 'd14;
assign strg_ub_tb_read_addr_gen_0_strides[0] = 'd1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[0] = 'd1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[1] = 'd4;
assign strg_ub_loops_buf2out_read_0_ranges[1] = 'd4;
assign strg_ub_tb_read_addr_gen_0_strides[1] = 'd1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[1] = 'd1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[2] = 'd-1;
assign strg_ub_loops_buf2out_read_0_ranges[2] = 'd-1;
assign strg_ub_tb_read_addr_gen_0_strides[2] = 'd-95;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[2] = 'd-95;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[0] = 'd14;
assign strg_ub_loops_buf2out_read_1_ranges[0] = 'd14;
assign strg_ub_tb_read_addr_gen_1_strides[0] = 'd1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[0] = 'd1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[1] = 'd4;
assign strg_ub_loops_buf2out_read_1_ranges[1] = 'd4;
assign strg_ub_tb_read_addr_gen_1_strides[1] = 'd1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[1] = 'd1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[2] = 'd-1;
assign strg_ub_loops_buf2out_read_1_ranges[2] = 'd-1;
assign strg_ub_tb_read_addr_gen_1_strides[2] = 'd-95;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[2] = 'd-95;

assign strg_ub_agg_read_addr_gen_0_starting_addr = 'b0;
assign strg_ub_input_addr_gen_starting_addr = 'b0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr = 'b100;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality = 'b11;
assign strg_ub_loops_in2buf_autovec_write_dimensionality = 'b11;
assign strg_ub_output_addr_gen_starting_addr = 'b0;
assign strg_ub_tb_write_addr_gen_0_starting_addr = 'b0;
assign strg_ub_tb_write_addr_gen_1_starting_addr = 'b0;
assign strg_ub_out_port_sel_addr_starting_addr = 'b0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr = 'b11101;
assign loops_buf2out_autovec_read_dimensionality = 'b100;
assign strg_ub_loops_buf2out_out_sel_dimensionality = 'b100;
assign strg_ub_agg_write_addr_gen_0_starting_addr = 'b0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr = 'b0;
assign strg_ub_loops_in2buf_0_dimensionality = 'b11;
assign strg_ub_tb_read_addr_gen_0_starting_addr = 'b0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr = 'b100000;
assign strg_ub_loops_buf2out_read_0_dimensionality = 'b11;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality = 'b11;
assign strg_ub_tb_read_addr_gen_1_starting_addr = 'b10000;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr = 'b100000;
assign strg_ub_loops_buf2out_read_1_dimensionality = 'b11;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality = 'b11;
assign chain_idx_input = 'b0;
assign chain_idx_output = 'b0;
assign enable_chain_input = 'b0;
assign enable_chain_output = 'b0;
assign chain_valid_in_reg_sel = 'b1;
assign chain_valid_in_reg_value = 'b0;
assign flush_reg_sel = 'b1;
assign flush_reg_value = 'b0;
assign ren_in_reg_sel = 'b1;
assign ren_in_reg_value = 'b0;
assign wen_in_reg_sel = 'b1;
assign wen_in_reg_value = 'b0;
assign mode = 'b0;
assign tile_en = 'b1;
assign strg_ub_loops_in2buf_0_ranges[0] = 'b10;
assign strg_ub_agg_write_addr_gen_0_strides[0] = 'b1;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[0] = 'b1;
assign strg_ub_loops_in2buf_0_ranges[1] = 'b11110;
assign strg_ub_agg_write_addr_gen_0_strides[1] = '0b11;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[1] = 'b1;
assign strg_ub_loops_in2buf_0_ranges[2] = '0b1;
assign strg_ub_agg_write_addr_gen_0_strides[2] = '0b11;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[2] = '0b1111111;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[0] = 'b10;
assign strg_ub_agg_read_addr_gen_0_strides[0] = 'b100;
assign strg_ub_loops_in2buf_autovec_write_ranges[0] = 'b10;
assign strg_ub_input_addr_gen_strides[0] = 'b1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[0] = 'b100;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[1] = 'b110;
assign strg_ub_agg_read_addr_gen_0_strides[1] = 'b100;
assign strg_ub_loops_in2buf_autovec_write_ranges[1] = 'b110;
assign strg_ub_input_addr_gen_strides[1] = 'b1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[1] = 'b100;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[2] = '0b1;
assign strg_ub_agg_read_addr_gen_0_strides[2] = '0b1111100;
assign strg_ub_loops_in2buf_autovec_write_ranges[2] = '0b1;
assign strg_ub_input_addr_gen_strides[2] = '0b11111;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[2] = '0b1111100;
assign strg_ub_loops_buf2out_autovec_read_ranges[0] = 'b0;
assign strg_ub_output_addr_gen_strides[0] = 'b100;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[0] = 'b10;
assign strg_ub_loops_buf2out_out_sel_ranges[0] = 'b0;
assign strg_ub_out_port_sel_addr_strides[0] = 'b1;
assign strg_ub_tb_write_addr_gen_0_strides[0] = 'b1;
assign strg_ub_tb_write_addr_gen_1_strides[0] = 'b1;
assign strg_ub_loops_buf2out_autovec_read_ranges[1] = 'b10;
assign strg_ub_output_addr_gen_strides[1] = '0b11;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[1] = 'b10;
assign strg_ub_loops_buf2out_out_sel_ranges[1] = 'b10;
assign strg_ub_out_port_sel_addr_strides[1] = '0b1;
assign strg_ub_tb_write_addr_gen_0_strides[1] = '0b1;
assign strg_ub_tb_write_addr_gen_1_strides[1] = '0b1;
assign strg_ub_loops_buf2out_autovec_read_ranges[2] = 'b100;
assign strg_ub_output_addr_gen_strides[2] = '0b11;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[2] = 'b10;
assign strg_ub_loops_buf2out_out_sel_ranges[2] = 'b100;
assign strg_ub_out_port_sel_addr_strides[2] = '0b1;
assign strg_ub_tb_write_addr_gen_0_strides[2] = '0b1;
assign strg_ub_tb_write_addr_gen_1_strides[2] = '0b1;
assign strg_ub_loops_buf2out_autovec_read_ranges[3] = '0b1;
assign strg_ub_output_addr_gen_strides[3] = '0b11011;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[3] = '0b1011110;
assign strg_ub_loops_buf2out_out_sel_ranges[3] = '0b1;
assign strg_ub_out_port_sel_addr_strides[3] = '0b1;
assign strg_ub_tb_write_addr_gen_0_strides[3] = '0b1;
assign strg_ub_tb_write_addr_gen_1_strides[3] = '0b1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[0] = 'b1110;
assign strg_ub_loops_buf2out_read_0_ranges[0] = 'b1110;
assign strg_ub_tb_read_addr_gen_0_strides[0] = 'b1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[0] = 'b1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[1] = 'b100;
assign strg_ub_loops_buf2out_read_0_ranges[1] = 'b100;
assign strg_ub_tb_read_addr_gen_0_strides[1] = 'b1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[1] = 'b1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[2] = '0b1;
assign strg_ub_loops_buf2out_read_0_ranges[2] = '0b1;
assign strg_ub_tb_read_addr_gen_0_strides[2] = '0b1011111;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[2] = '0b1011111;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[0] = 'b1110;
assign strg_ub_loops_buf2out_read_1_ranges[0] = 'b1110;
assign strg_ub_tb_read_addr_gen_1_strides[0] = 'b1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[0] = 'b1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[1] = 'b100;
assign strg_ub_loops_buf2out_read_1_ranges[1] = 'b100;
assign strg_ub_tb_read_addr_gen_1_strides[1] = 'b1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[1] = 'b1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[2] = '0b1;
assign strg_ub_loops_buf2out_read_1_ranges[2] = '0b1;
assign strg_ub_tb_read_addr_gen_1_strides[2] = '0b1011111;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[2] = '0b1011111;

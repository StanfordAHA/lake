assign strg_ub_agg_read_addr_gen_0_starting_addr = 8'b0;
assign strg_ub_input_addr_gen_starting_addr = 16'b0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr = 16'b100;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality = 3'b11;
assign strg_ub_loops_in2buf_autovec_write_dimensionality = 4'b11;
assign strg_ub_output_addr_gen_starting_addr = 16'b0;
assign strg_ub_tb_write_addr_gen_0_starting_addr = 6'b0;
assign strg_ub_tb_write_addr_gen_1_starting_addr = 6'b0;
assign strg_ub_out_port_sel_addr_starting_addr = 1'b0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr = 16'b11101;
assign strg_ub_loops_buf2out_autovec_read_dimensionality = 4'b100;
assign strg_ub_loops_buf2out_out_sel_dimensionality = 2'b100;
assign strg_ub_agg_write_addr_gen_0_starting_addr = 4'b0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr = 4'b0;
assign strg_ub_loops_in2buf_0_dimensionality = 3'b11;
assign strg_ub_tb_read_addr_gen_0_starting_addr = 6'b0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr = 16'b100000;
assign strg_ub_loops_buf2out_read_0_dimensionality = 2'b11;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality = 2'b11;
assign strg_ub_tb_read_addr_gen_1_starting_addr = 6'b10000;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr = 16'b100000;
assign strg_ub_loops_buf2out_read_1_dimensionality = 2'b11;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality = 2'b11;
assign mode = 2'b0;
assign tile_en = 1'b1;
assign strg_ub_loops_in2buf_0_ranges[0] = 4'b10;
assign strg_ub_agg_write_addr_gen_0_strides[0] = 4'b1;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[0] = 4'b1;
assign strg_ub_loops_in2buf_0_ranges[1] = 4'b11110;
assign strg_ub_agg_write_addr_gen_0_strides[1] = 4'b11;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[1] = 4'b1;
assign strg_ub_loops_in2buf_0_ranges[2] = 4'b1;
assign strg_ub_agg_write_addr_gen_0_strides[2] = 4'b11;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides[2] = 4'b1111111;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[0] = 8'b10;
assign strg_ub_agg_read_addr_gen_0_strides[0] = 8'b100;
assign strg_ub_loops_in2buf_autovec_write_ranges[0] = 16'b10;
assign strg_ub_input_addr_gen_strides[0] = 16'b1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[0] = 16'b100;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[1] = 8'b110;
assign strg_ub_agg_read_addr_gen_0_strides[1] = 8'b100;
assign strg_ub_loops_in2buf_autovec_write_ranges[1] = 16'b110;
assign strg_ub_input_addr_gen_strides[1] = 16'b1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[1] = 16'b100;
assign strg_ub_loops_in2buf_autovec_read_0_ranges[2] = 8'b1;
assign strg_ub_agg_read_addr_gen_0_strides[2] = 8'b1111100;
assign strg_ub_loops_in2buf_autovec_write_ranges[2] = 16'b1;
assign strg_ub_input_addr_gen_strides[2] = 16'b11111;
assign strg_ub_input_sched_gen_sched_addr_gen_strides[2] = 16'b1111100;
assign strg_ub_loops_buf2out_autovec_read_ranges[0] = 16'b0;
assign strg_ub_output_addr_gen_strides[0] = 16'b100;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[0] = 16'b10;
assign strg_ub_loops_buf2out_out_sel_ranges[0] = 1'b0;
assign strg_ub_out_port_sel_addr_strides[0] = 1'b1;
assign strg_ub_tb_write_addr_gen_0_strides[0] = 6'b1;
assign strg_ub_tb_write_addr_gen_1_strides[0] = 6'b1;
assign strg_ub_loops_buf2out_autovec_read_ranges[1] = 16'b10;
assign strg_ub_output_addr_gen_strides[1] = 16'b11;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[1] = 16'b10;
assign strg_ub_loops_buf2out_out_sel_ranges[1] = 1'b10;
assign strg_ub_out_port_sel_addr_strides[1] = 1'b1;
assign strg_ub_tb_write_addr_gen_0_strides[1] = 6'b1;
assign strg_ub_tb_write_addr_gen_1_strides[1] = 6'b1;
assign strg_ub_loops_buf2out_autovec_read_ranges[2] = 16'b100;
assign strg_ub_output_addr_gen_strides[2] = 16'b11;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[2] = 16'b10;
assign strg_ub_loops_buf2out_out_sel_ranges[2] = 1'b100;
assign strg_ub_out_port_sel_addr_strides[2] = 1'b1;
assign strg_ub_tb_write_addr_gen_0_strides[2] = 6'b1;
assign strg_ub_tb_write_addr_gen_1_strides[2] = 6'b1;
assign strg_ub_loops_buf2out_autovec_read_ranges[3] = 16'b1;
assign strg_ub_output_addr_gen_strides[3] = 16'b11011;
assign strg_ub_output_sched_gen_sched_addr_gen_strides[3] = 16'b1011110;
assign strg_ub_loops_buf2out_out_sel_ranges[3] = 1'b1;
assign strg_ub_out_port_sel_addr_strides[3] = 1'b1;
assign strg_ub_tb_write_addr_gen_0_strides[3] = 6'b1;
assign strg_ub_tb_write_addr_gen_1_strides[3] = 6'b1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[0] = 6'b1110;
assign strg_ub_loops_buf2out_read_0_ranges[0] = 16'b1110;
assign strg_ub_tb_read_addr_gen_0_strides[0] = 6'b1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[0] = 16'b1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[1] = 6'b100;
assign strg_ub_loops_buf2out_read_0_ranges[1] = 16'b100;
assign strg_ub_tb_read_addr_gen_0_strides[1] = 6'b1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[1] = 16'b1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges[2] = 6'b1;
assign strg_ub_loops_buf2out_read_0_ranges[2] = 16'b1;
assign strg_ub_tb_read_addr_gen_0_strides[2] = 6'b1011111;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides[2] = 16'b1011111;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[0] = 6'b1110;
assign strg_ub_loops_buf2out_read_1_ranges[0] = 16'b1110;
assign strg_ub_tb_read_addr_gen_1_strides[0] = 6'b1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[0] = 16'b1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[1] = 6'b100;
assign strg_ub_loops_buf2out_read_1_ranges[1] = 16'b100;
assign strg_ub_tb_read_addr_gen_1_strides[1] = 6'b1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[1] = 16'b1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges[2] = 6'b1;
assign strg_ub_loops_buf2out_read_1_ranges[2] = 16'b1;
assign strg_ub_tb_read_addr_gen_1_strides[2] = 6'b1011111;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides[2] = 16'b1011111;

wire [15:0] strg_ub_agg_read_addr_gen_0_starting_addr = 0;
wire [15:0] strg_ub_input_addr_gen_starting_addr = 0;
wire [15:0] strg_ub_input_sched_gen_sched_addr_gen_starting_addr = 4;
wire [3:0] strg_ub_loops_in2buf_autovec_read_0_dimensionality = 3;
wire [3:0] strg_ub_loops_in2buf_autovec_write_dimensionality = 3;
wire [15:0] strg_ub_output_addr_gen_starting_addr = 0;
wire [15:0] strg_ub_tb_write_addr_gen_0_starting_addr = 0;
wire [15:0] strg_ub_tb_write_addr_gen_1_starting_addr = 0;
wire [15:0] strg_ub_out_port_sel_addr_starting_addr = 0;
wire [15:0] strg_ub_output_sched_gen_sched_addr_gen_starting_addr = 29;
wire [3:0] strg_ub_loops_buf2out_autovec_read_dimensionality = 4;
wire [3:0] strg_ub_loops_buf2out_out_sel_dimensionality = 4;
wire [15:0] strg_ub_agg_write_addr_gen_0_starting_addr = 0;
wire [15:0] strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr = 0;
wire [3:0] strg_ub_loops_in2buf_0_dimensionality = 4;
wire [15:0] strg_ub_tb_read_addr_gen_0_starting_addr = 0;
wire [15:0] strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr = 33;
wire [3:0] strg_ub_loops_buf2out_read_0_dimensionality = 4;
wire [3:0] strg_ub_loops_buf2out_autovec_write_0_dimensionality = 4;
wire [15:0] strg_ub_tb_read_addr_gen_1_starting_addr = 0;
wire [15:0] strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr = 33;
wire [3:0] strg_ub_loops_buf2out_read_1_dimensionality = 4;
wire [3:0] strg_ub_loops_buf2out_autovec_write_1_dimensionality = 4;
wire [1:0] mode = 0;
wire [0:0] tile_en = 1;
wire [15:0] strg_ub_loops_in2buf_0_ranges_0 = 2;
wire [15:0] strg_ub_agg_write_addr_gen_0_strides_0 = 1;
wire [15:0] strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_0 = 1;
wire [15:0] strg_ub_loops_in2buf_0_ranges_1 = 2;
wire [15:0] strg_ub_agg_write_addr_gen_0_strides_1 = -3;
wire [15:0] strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_1 = 1;
wire [15:0] strg_ub_loops_in2buf_0_ranges_2 = 6;
wire [15:0] strg_ub_agg_write_addr_gen_0_strides_2 = -3;
wire [15:0] strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_2 = 1;
wire [15:0] strg_ub_loops_in2buf_0_ranges_3 = -1;
wire [15:0] strg_ub_agg_write_addr_gen_0_strides_3 = -3;
wire [15:0] strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_3 = -127;
wire [15:0] strg_ub_loops_in2buf_autovec_read_0_ranges_0 = 2;
wire [15:0] strg_ub_agg_read_addr_gen_0_strides_0 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_write_ranges_0 = 2;
wire [15:0] strg_ub_input_addr_gen_strides_0 = 1;
wire [15:0] strg_ub_input_sched_gen_sched_addr_gen_strides_0 = 4;
wire [15:0] strg_ub_loops_in2buf_autovec_read_0_ranges_1 = 6;
wire [15:0] strg_ub_agg_read_addr_gen_0_strides_1 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_write_ranges_1 = 6;
wire [15:0] strg_ub_input_addr_gen_strides_1 = 1;
wire [15:0] strg_ub_input_sched_gen_sched_addr_gen_strides_1 = 4;
wire [15:0] strg_ub_loops_in2buf_autovec_read_0_ranges_2 = -1;
wire [15:0] strg_ub_agg_read_addr_gen_0_strides_2 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_write_ranges_2 = -1;
wire [15:0] strg_ub_input_addr_gen_strides_2 = -31;
wire [15:0] strg_ub_input_sched_gen_sched_addr_gen_strides_2 = -124;
wire [15:0] strg_ub_loops_buf2out_autovec_read_ranges_0 = 0;
wire [15:0] strg_ub_output_addr_gen_strides_0 = 4;
wire [15:0] strg_ub_output_sched_gen_sched_addr_gen_strides_0 = 2;
wire [15:0] strg_ub_loops_buf2out_out_sel_ranges_0 = 0;
wire [15:0] strg_ub_out_port_sel_addr_strides_0 = 1;
wire [15:0] strg_ub_tb_write_addr_gen_0_strides_0 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_write_0_ranges_0 = 0;
wire [15:0] strg_ub_tb_write_addr_gen_1_strides_0 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_write_1_ranges_0 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_read_ranges_1 = 2;
wire [15:0] strg_ub_output_addr_gen_strides_1 = -3;
wire [15:0] strg_ub_output_sched_gen_sched_addr_gen_strides_1 = 2;
wire [15:0] strg_ub_loops_buf2out_out_sel_ranges_1 = 2;
wire [15:0] strg_ub_out_port_sel_addr_strides_1 = -1;
wire [15:0] strg_ub_tb_write_addr_gen_0_strides_1 = 1;
wire [15:0] strg_ub_loops_buf2out_autovec_write_0_ranges_1 = 2;
wire [15:0] strg_ub_tb_write_addr_gen_1_strides_1 = 1;
wire [15:0] strg_ub_loops_buf2out_autovec_write_1_ranges_1 = 2;
wire [15:0] strg_ub_loops_buf2out_autovec_read_ranges_2 = 4;
wire [15:0] strg_ub_output_addr_gen_strides_2 = -3;
wire [15:0] strg_ub_output_sched_gen_sched_addr_gen_strides_2 = 2;
wire [15:0] strg_ub_loops_buf2out_out_sel_ranges_2 = 4;
wire [15:0] strg_ub_out_port_sel_addr_strides_2 = -1;
wire [15:0] strg_ub_tb_write_addr_gen_0_strides_2 = -3;
wire [15:0] strg_ub_loops_buf2out_autovec_write_0_ranges_2 = 4;
wire [15:0] strg_ub_tb_write_addr_gen_1_strides_2 = -3;
wire [15:0] strg_ub_loops_buf2out_autovec_write_1_ranges_2 = 4;
wire [15:0] strg_ub_loops_buf2out_autovec_read_ranges_3 = -1;
wire [15:0] strg_ub_output_addr_gen_strides_3 = -27;
wire [15:0] strg_ub_output_sched_gen_sched_addr_gen_strides_3 = -94;
wire [15:0] strg_ub_loops_buf2out_out_sel_ranges_3 = -1;
wire [15:0] strg_ub_out_port_sel_addr_strides_3 = -1;
wire [15:0] strg_ub_tb_write_addr_gen_0_strides_3 = -3;
wire [15:0] strg_ub_loops_buf2out_autovec_write_0_ranges_3 = -1;
wire [15:0] strg_ub_tb_write_addr_gen_1_strides_3 = -3;
wire [15:0] strg_ub_loops_buf2out_autovec_write_1_ranges_3 = -1;
wire [15:0] strg_ub_loops_buf2out_read_0_ranges_0 = 2;
wire [15:0] strg_ub_tb_read_addr_gen_0_strides_0 = 1;
wire [15:0] strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_0 = 1;
wire [15:0] strg_ub_loops_buf2out_read_0_ranges_1 = 2;
wire [15:0] strg_ub_tb_read_addr_gen_0_strides_1 = 1;
wire [15:0] strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_1 = 1;
wire [15:0] strg_ub_loops_buf2out_read_0_ranges_2 = 4;
wire [15:0] strg_ub_tb_read_addr_gen_0_strides_2 = -15;
wire [15:0] strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_2 = 1;
wire [15:0] strg_ub_loops_buf2out_read_0_ranges_3 = -1;
wire [15:0] strg_ub_tb_read_addr_gen_0_strides_3 = -15;
wire [15:0] strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_3 = -95;
wire [15:0] strg_ub_loops_buf2out_read_1_ranges_0 = 2;
wire [15:0] strg_ub_tb_read_addr_gen_1_strides_0 = 1;
wire [15:0] strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_0 = 1;
wire [15:0] strg_ub_loops_buf2out_read_1_ranges_1 = 2;
wire [15:0] strg_ub_tb_read_addr_gen_1_strides_1 = 1;
wire [15:0] strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_1 = 1;
wire [15:0] strg_ub_loops_buf2out_read_1_ranges_2 = 4;
wire [15:0] strg_ub_tb_read_addr_gen_1_strides_2 = -15;
wire [15:0] strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_2 = 1;
wire [15:0] strg_ub_loops_buf2out_read_1_ranges_3 = -1;
wire [15:0] strg_ub_tb_read_addr_gen_1_strides_3 = -15;
wire [15:0] strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_3 = -95;
wire [15:0] strg_ub_loops_buf2out_autovec_write_1_ranges_4 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_write_1_ranges_5 = 0;
wire [15:0] strg_ub_input_addr_gen_strides_3 = 0;
wire [15:0] strg_ub_input_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_input_addr_gen_strides_5 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_0_strides_4 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_0_strides_5 = 0;
wire [15:0] strg_ub_loops_buf2out_read_1_ranges_4 = 0;
wire [15:0] strg_ub_loops_buf2out_read_1_ranges_5 = 0;
wire [15:0] strg_ub_out_port_sel_addr_strides_4 = 0;
wire [15:0] strg_ub_out_port_sel_addr_strides_5 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_0_ranges_3 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_0_ranges_4 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_0_ranges_5 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_write_0_ranges_4 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_write_0_ranges_5 = 0;
wire [15:0] strg_ub_input_sched_gen_sched_addr_gen_strides_3 = 0;
wire [15:0] strg_ub_input_sched_gen_sched_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_input_sched_gen_sched_addr_gen_strides_5 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_0 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_1 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_2 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_3 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_5 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_1_ranges_0 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_1_ranges_1 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_1_ranges_2 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_1_ranges_3 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_1_ranges_4 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_1_ranges_5 = 0;
wire [15:0] strg_ub_port_sel_addr_starting_addr = 0;
wire [15:0] strg_ub_agg_read_addr_gen_0_strides_3 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_0_strides_4 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_0_strides_5 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_1_starting_addr = 0;
wire [15:0] strg_ub_tb_write_addr_gen_0_strides_4 = 0;
wire [15:0] strg_ub_tb_write_addr_gen_0_strides_5 = 0;
wire [15:0] strg_ub_loops_buf2out_out_sel_ranges_4 = 0;
wire [15:0] strg_ub_loops_buf2out_out_sel_ranges_5 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_write_ranges_3 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_write_ranges_4 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_write_ranges_5 = 0;
wire [15:0] strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_5 = 0;
wire [15:0] strg_ub_loops_in2buf_0_ranges_4 = 0;
wire [15:0] strg_ub_loops_in2buf_0_ranges_5 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_1_strides_0 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_1_strides_1 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_1_strides_2 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_1_strides_3 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_1_strides_4 = 0;
wire [15:0] strg_ub_agg_read_addr_gen_1_strides_5 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_1_starting_addr = 0;
wire [15:0] strg_ub_tb_write_addr_gen_1_strides_4 = 0;
wire [15:0] strg_ub_tb_write_addr_gen_1_strides_5 = 0;
wire [15:0] strg_ub_tb_read_addr_gen_0_strides_4 = 0;
wire [15:0] strg_ub_tb_read_addr_gen_0_strides_5 = 0;
wire [15:0] strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_5 = 0;
wire [15:0] strg_ub_loops_in2buf_autovec_read_1_dimensionality = 0;
wire [15:0] strg_ub_port_sel_addr_strides_0 = 0;
wire [15:0] strg_ub_port_sel_addr_strides_1 = 0;
wire [15:0] strg_ub_port_sel_addr_strides_2 = 0;
wire [15:0] strg_ub_port_sel_addr_strides_3 = 0;
wire [15:0] strg_ub_port_sel_addr_strides_4 = 0;
wire [15:0] strg_ub_port_sel_addr_strides_5 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_read_ranges_4 = 0;
wire [15:0] strg_ub_loops_buf2out_autovec_read_ranges_5 = 0;
wire [15:0] strg_ub_loops_in2buf_1_dimensionality = 0;
wire [15:0] strg_ub_loops_buf2out_read_0_ranges_4 = 0;
wire [15:0] strg_ub_loops_buf2out_read_0_ranges_5 = 0;
wire [15:0] strg_ub_tb_read_addr_gen_1_strides_4 = 0;
wire [15:0] strg_ub_tb_read_addr_gen_1_strides_5 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_1_sched_addr_gen_starting_addr = 0;
wire [15:0] strg_ub_agg_write_addr_gen_1_strides_0 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_1_strides_1 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_1_strides_2 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_1_strides_3 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_1_strides_4 = 0;
wire [15:0] strg_ub_agg_write_addr_gen_1_strides_5 = 0;
wire [15:0] strg_ub_output_sched_gen_sched_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_output_sched_gen_sched_addr_gen_strides_5 = 0;
wire [15:0] strg_ub_output_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_output_addr_gen_strides_5 = 0;
wire [15:0] strg_ub_loops_in2buf_1_ranges_0 = 0;
wire [15:0] strg_ub_loops_in2buf_1_ranges_1 = 0;
wire [15:0] strg_ub_loops_in2buf_1_ranges_2 = 0;
wire [15:0] strg_ub_loops_in2buf_1_ranges_3 = 0;
wire [15:0] strg_ub_loops_in2buf_1_ranges_4 = 0;
wire [15:0] strg_ub_loops_in2buf_1_ranges_5 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_4 = 0;
wire [15:0] strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_5 = 0;

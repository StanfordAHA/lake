assign strg_ub_agg_read_addr_gen_0_starting_addr = 8'h0;
assign strg_ub_input_addr_gen_starting_addr = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr = 16'h4;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality = 3'h3;
assign strg_ub_loops_in2buf_autovec_write_dimensionality = 4'h3;
assign strg_ub_output_addr_gen_starting_addr = 16'h0;
assign strg_ub_tb_write_addr_gen_0_starting_addr = 6'h0;
assign strg_ub_tb_write_addr_gen_1_starting_addr = 6'h0;
assign strg_ub_out_port_sel_addr_starting_addr = 1'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr = 16'h1D;
assign strg_ub_loops_buf2out_autovec_read_dimensionality = 4'h4;
assign strg_ub_loops_buf2out_out_sel_dimensionality = 2'h4;
assign strg_ub_agg_write_addr_gen_0_starting_addr = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr = 4'h0;
assign strg_ub_loops_in2buf_0_dimensionality = 3'h3;
assign strg_ub_tb_read_addr_gen_0_starting_addr = 6'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr = 16'h20;
assign strg_ub_loops_buf2out_read_0_dimensionality = 2'h3;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality = 2'h3;
assign strg_ub_tb_read_addr_gen_1_starting_addr = 6'h10;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr = 16'h20;
assign strg_ub_loops_buf2out_read_1_dimensionality = 2'h3;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality = 2'h3;
assign mode = 2'h0;
assign tile_en = 1'h1;
assign strg_ub_loops_in2buf_0_ranges_0 = 4'h2;
assign strg_ub_agg_write_addr_gen_0_strides_0 = 4'h1;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_0 = 4'h1;
assign strg_ub_loops_in2buf_0_ranges_1 = 4'hE;
assign strg_ub_agg_write_addr_gen_0_strides_1 = 4'h3;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_1 = 4'h1;
assign strg_ub_loops_in2buf_0_ranges_2 = 4'h1;
assign strg_ub_agg_write_addr_gen_0_strides_2 = 4'h3;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_2 = 4'h1;
assign strg_ub_loops_in2buf_autovec_read_0_ranges_0 = 8'h2;
assign strg_ub_agg_read_addr_gen_0_strides_0 = 8'h4;
assign strg_ub_loops_in2buf_autovec_write_ranges_0 = 16'h2;
assign strg_ub_input_addr_gen_strides_0 = 16'h1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides_0 = 16'h4;
assign strg_ub_loops_in2buf_autovec_read_0_ranges_1 = 8'h6;
assign strg_ub_agg_read_addr_gen_0_strides_1 = 8'h4;
assign strg_ub_loops_in2buf_autovec_write_ranges_1 = 16'h6;
assign strg_ub_input_addr_gen_strides_1 = 16'h1;
assign strg_ub_input_sched_gen_sched_addr_gen_strides_1 = 16'h4;
assign strg_ub_loops_in2buf_autovec_read_0_ranges_2 = 8'h1;
assign strg_ub_agg_read_addr_gen_0_strides_2 = 8'h7C;
assign strg_ub_loops_in2buf_autovec_write_ranges_2 = 16'h1;
assign strg_ub_input_addr_gen_strides_2 = 16'h1F;
assign strg_ub_input_sched_gen_sched_addr_gen_strides_2 = 16'h7C;
assign strg_ub_loops_buf2out_autovec_read_ranges_0 = 16'h0;
assign strg_ub_output_addr_gen_strides_0 = 16'h4;
assign strg_ub_output_sched_gen_sched_addr_gen_strides_0 = 16'h2;
assign strg_ub_loops_buf2out_out_sel_ranges_0 = 1'h0;
assign strg_ub_out_port_sel_addr_strides_0 = 1'h1;
assign strg_ub_tb_write_addr_gen_0_strides_0 = 6'h1;
assign strg_ub_tb_write_addr_gen_1_strides_0 = 6'h1;
assign strg_ub_loops_buf2out_autovec_read_ranges_1 = 16'h2;
assign strg_ub_output_addr_gen_strides_1 = 16'h3;
assign strg_ub_output_sched_gen_sched_addr_gen_strides_1 = 16'h2;
assign strg_ub_loops_buf2out_out_sel_ranges_1 = 1'h2;
assign strg_ub_out_port_sel_addr_strides_1 = 1'h1;
assign strg_ub_tb_write_addr_gen_0_strides_1 = 6'h1;
assign strg_ub_tb_write_addr_gen_1_strides_1 = 6'h1;
assign strg_ub_loops_buf2out_autovec_read_ranges_2 = 16'h4;
assign strg_ub_output_addr_gen_strides_2 = 16'h3;
assign strg_ub_output_sched_gen_sched_addr_gen_strides_2 = 16'h2;
assign strg_ub_loops_buf2out_out_sel_ranges_2 = 1'h4;
assign strg_ub_out_port_sel_addr_strides_2 = 1'h1;
assign strg_ub_tb_write_addr_gen_0_strides_2 = 6'h1;
assign strg_ub_tb_write_addr_gen_1_strides_2 = 6'h1;
assign strg_ub_loops_buf2out_autovec_read_ranges_3 = 16'h1;
assign strg_ub_output_addr_gen_strides_3 = 16'h1B;
assign strg_ub_output_sched_gen_sched_addr_gen_strides_3 = 16'h5E;
assign strg_ub_loops_buf2out_out_sel_ranges_3 = 1'h1;
assign strg_ub_out_port_sel_addr_strides_3 = 1'h1;
assign strg_ub_tb_write_addr_gen_0_strides_3 = 6'h1;
assign strg_ub_tb_write_addr_gen_1_strides_3 = 6'h1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges_0 = 6'hE;
assign strg_ub_loops_buf2out_read_0_ranges_0 = 16'hE;
assign strg_ub_tb_read_addr_gen_0_strides_0 = 6'h1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_0 = 16'h1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges_1 = 6'h4;
assign strg_ub_loops_buf2out_read_0_ranges_1 = 16'h4;
assign strg_ub_tb_read_addr_gen_0_strides_1 = 6'h1;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_1 = 16'h1;
assign strg_ub_loops_buf2out_autovec_write_0_ranges_2 = 6'h1;
assign strg_ub_loops_buf2out_read_0_ranges_2 = 16'h1;
assign strg_ub_tb_read_addr_gen_0_strides_2 = 6'h5F;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_2 = 16'h5F;
assign strg_ub_loops_buf2out_autovec_write_1_ranges_0 = 6'hE;
assign strg_ub_loops_buf2out_read_1_ranges_0 = 16'hE;
assign strg_ub_tb_read_addr_gen_1_strides_0 = 6'h1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_0 = 16'h1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges_1 = 6'h4;
assign strg_ub_loops_buf2out_read_1_ranges_1 = 16'h4;
assign strg_ub_tb_read_addr_gen_1_strides_1 = 6'h1;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_1 = 16'h1;
assign strg_ub_loops_buf2out_autovec_write_1_ranges_2 = 6'h1;
assign strg_ub_loops_buf2out_read_1_ranges_2 = 16'h1;
assign strg_ub_tb_read_addr_gen_1_strides_2 = 6'h5F;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_2 = 16'h5F;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality_0 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality_1 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality_2 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality_3 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality_4 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_0_dimensionality_5 = 2'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr_0 = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr_1 = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr_2 = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr_3 = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr_4 = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_starting_addr_5 = 16'h0;
assign strg_ub_agg_read_addr_gen_0_starting_addr_0 = 8'h0;
assign strg_ub_agg_read_addr_gen_0_starting_addr_1 = 8'h0;
assign strg_ub_agg_read_addr_gen_0_starting_addr_2 = 8'h0;
assign strg_ub_agg_read_addr_gen_0_starting_addr_3 = 8'h0;
assign strg_ub_agg_read_addr_gen_0_starting_addr_4 = 8'h0;
assign strg_ub_agg_read_addr_gen_0_starting_addr_5 = 8'h0;
assign strg_ub_loops_buf2out_read_1_ranges_3 = 16'h0;
assign strg_ub_loops_buf2out_read_1_ranges_4 = 16'h0;
assign strg_ub_loops_buf2out_read_1_ranges_5 = 16'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_0 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_1 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_2 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_3 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_4 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_strides_5 = 4'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_3 = 16'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_4 = 16'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_strides_5 = 16'h0;
assign strg_ub_tb_read_addr_gen_1_strides_3 = 6'h0;
assign strg_ub_tb_read_addr_gen_1_strides_4 = 6'h0;
assign strg_ub_tb_read_addr_gen_1_strides_5 = 6'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr_0 = 16'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr_1 = 16'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr_2 = 16'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr_3 = 16'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr_4 = 16'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_starting_addr_5 = 16'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_strides_4 = 16'h0;
assign strg_ub_output_sched_gen_sched_addr_gen_strides_5 = 16'h0;
assign strg_ub_loops_in2buf_0_dimensionality_0 = 3'h0;
assign strg_ub_loops_in2buf_0_dimensionality_1 = 3'h0;
assign strg_ub_loops_in2buf_0_dimensionality_2 = 3'h0;
assign strg_ub_loops_in2buf_0_dimensionality_3 = 3'h0;
assign strg_ub_loops_in2buf_0_dimensionality_4 = 3'h0;
assign strg_ub_loops_in2buf_0_dimensionality_5 = 3'h0;
assign strg_ub_loops_buf2out_autovec_write_1_ranges_3 = 6'h0;
assign strg_ub_loops_buf2out_autovec_write_1_ranges_4 = 6'h0;
assign strg_ub_loops_buf2out_autovec_write_1_ranges_5 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_strides_3 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_strides_4 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_strides_5 = 6'h0;
assign strg_ub_agg_write_addr_gen_1_starting_addr_0 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_starting_addr_1 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_starting_addr_2 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_starting_addr_3 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_starting_addr_4 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_starting_addr_5 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr_0 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr_1 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr_2 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr_3 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr_4 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_starting_addr_5 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_3 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_4 = 4'h0;
assign strg_ub_agg_write_sched_gen_0_sched_addr_gen_strides_5 = 4'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_strides_3 = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_strides_4 = 16'h0;
assign strg_ub_input_sched_gen_sched_addr_gen_strides_5 = 16'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_starting_addr_0 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_starting_addr_1 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_starting_addr_2 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_starting_addr_3 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_starting_addr_4 = 4'h0;
assign strg_ub_agg_write_sched_gen_1_sched_addr_gen_starting_addr_5 = 4'h0;
assign strg_ub_loops_buf2out_autovec_write_0_ranges_3 = 6'h0;
assign strg_ub_loops_buf2out_autovec_write_0_ranges_4 = 6'h0;
assign strg_ub_loops_buf2out_autovec_write_0_ranges_5 = 6'h0;
assign strg_ub_loops_buf2out_read_0_ranges_3 = 16'h0;
assign strg_ub_loops_buf2out_read_0_ranges_4 = 16'h0;
assign strg_ub_loops_buf2out_read_0_ranges_5 = 16'h0;
assign strg_ub_loops_buf2out_autovec_read_ranges_4 = 16'h0;
assign strg_ub_loops_buf2out_autovec_read_ranges_5 = 16'h0;
assign strg_ub_loops_in2buf_autovec_write_ranges_3 = 16'h0;
assign strg_ub_loops_in2buf_autovec_write_ranges_4 = 16'h0;
assign strg_ub_loops_in2buf_autovec_write_ranges_5 = 16'h0;
assign strg_ub_loops_in2buf_autovec_read_0_ranges_3 = 8'h0;
assign strg_ub_loops_in2buf_autovec_read_0_ranges_4 = 8'h0;
assign strg_ub_loops_in2buf_autovec_read_0_ranges_5 = 8'h0;
assign strg_ub_tb_read_addr_gen_0_starting_addr_0 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_starting_addr_1 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_starting_addr_2 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_starting_addr_3 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_starting_addr_4 = 6'h0;
assign strg_ub_tb_read_addr_gen_0_starting_addr_5 = 6'h0;
assign strg_ub_out_port_sel_addr_strides_4 = 1'h0;
assign strg_ub_out_port_sel_addr_strides_5 = 1'h0;
assign strg_ub_loops_buf2out_autovec_read_dimensionality_0 = 4'h0;
assign strg_ub_loops_buf2out_autovec_read_dimensionality_1 = 4'h0;
assign strg_ub_loops_buf2out_autovec_read_dimensionality_2 = 4'h0;
assign strg_ub_loops_buf2out_autovec_read_dimensionality_3 = 4'h0;
assign strg_ub_loops_buf2out_autovec_read_dimensionality_4 = 4'h0;
assign strg_ub_loops_buf2out_autovec_read_dimensionality_5 = 4'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_3 = 16'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_4 = 16'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_strides_5 = 16'h0;
assign strg_ub_loops_buf2out_out_sel_ranges_4 = 1'h0;
assign strg_ub_loops_buf2out_out_sel_ranges_5 = 1'h0;
assign strg_ub_agg_read_addr_gen_1_starting_addr_0 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_starting_addr_1 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_starting_addr_2 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_starting_addr_3 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_starting_addr_4 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_starting_addr_5 = 8'h0;
assign strg_ub_agg_write_addr_gen_0_strides_3 = 4'h0;
assign strg_ub_agg_write_addr_gen_0_strides_4 = 4'h0;
assign strg_ub_agg_write_addr_gen_0_strides_5 = 4'h0;
assign strg_ub_loops_in2buf_autovec_read_1_dimensionality_0 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_1_dimensionality_1 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_1_dimensionality_2 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_1_dimensionality_3 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_1_dimensionality_4 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_1_dimensionality_5 = 3'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr_0 = 16'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr_1 = 16'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr_2 = 16'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr_3 = 16'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr_4 = 16'h0;
assign strg_ub_tb_read_sched_gen_0_sched_addr_gen_starting_addr_5 = 16'h0;
assign strg_ub_loops_buf2out_read_0_dimensionality_0 = 2'h0;
assign strg_ub_loops_buf2out_read_0_dimensionality_1 = 2'h0;
assign strg_ub_loops_buf2out_read_0_dimensionality_2 = 2'h0;
assign strg_ub_loops_buf2out_read_0_dimensionality_3 = 2'h0;
assign strg_ub_loops_buf2out_read_0_dimensionality_4 = 2'h0;
assign strg_ub_loops_buf2out_read_0_dimensionality_5 = 2'h0;
assign strg_ub_loops_buf2out_out_sel_dimensionality_0 = 2'h0;
assign strg_ub_loops_buf2out_out_sel_dimensionality_1 = 2'h0;
assign strg_ub_loops_buf2out_out_sel_dimensionality_2 = 2'h0;
assign strg_ub_loops_buf2out_out_sel_dimensionality_3 = 2'h0;
assign strg_ub_loops_buf2out_out_sel_dimensionality_4 = 2'h0;
assign strg_ub_loops_buf2out_out_sel_dimensionality_5 = 2'h0;
assign strg_ub_input_addr_gen_starting_addr_0 = 16'h0;
assign strg_ub_input_addr_gen_starting_addr_1 = 16'h0;
assign strg_ub_input_addr_gen_starting_addr_2 = 16'h0;
assign strg_ub_input_addr_gen_starting_addr_3 = 16'h0;
assign strg_ub_input_addr_gen_starting_addr_4 = 16'h0;
assign strg_ub_input_addr_gen_starting_addr_5 = 16'h0;
assign strg_ub_loops_in2buf_0_ranges_3 = 4'h0;
assign strg_ub_loops_in2buf_0_ranges_4 = 4'h0;
assign strg_ub_loops_in2buf_0_ranges_5 = 4'h0;
assign strg_ub_loops_in2buf_1_dimensionality_0 = 3'h0;
assign strg_ub_loops_in2buf_1_dimensionality_1 = 3'h0;
assign strg_ub_loops_in2buf_1_dimensionality_2 = 3'h0;
assign strg_ub_loops_in2buf_1_dimensionality_3 = 3'h0;
assign strg_ub_loops_in2buf_1_dimensionality_4 = 3'h0;
assign strg_ub_loops_in2buf_1_dimensionality_5 = 3'h0;
assign strg_ub_port_sel_addr_strides_0 = 1'h0;
assign strg_ub_port_sel_addr_strides_1 = 1'h0;
assign strg_ub_port_sel_addr_strides_2 = 1'h0;
assign strg_ub_port_sel_addr_strides_3 = 1'h0;
assign strg_ub_port_sel_addr_strides_4 = 1'h0;
assign strg_ub_port_sel_addr_strides_5 = 1'h0;
assign strg_ub_port_sel_addr_starting_addr_0 = 1'h0;
assign strg_ub_port_sel_addr_starting_addr_1 = 1'h0;
assign strg_ub_port_sel_addr_starting_addr_2 = 1'h0;
assign strg_ub_port_sel_addr_starting_addr_3 = 1'h0;
assign strg_ub_port_sel_addr_starting_addr_4 = 1'h0;
assign strg_ub_port_sel_addr_starting_addr_5 = 1'h0;
assign strg_ub_loops_in2buf_autovec_write_dimensionality_0 = 4'h0;
assign strg_ub_loops_in2buf_autovec_write_dimensionality_1 = 4'h0;
assign strg_ub_loops_in2buf_autovec_write_dimensionality_2 = 4'h0;
assign strg_ub_loops_in2buf_autovec_write_dimensionality_3 = 4'h0;
assign strg_ub_loops_in2buf_autovec_write_dimensionality_4 = 4'h0;
assign strg_ub_loops_in2buf_autovec_write_dimensionality_5 = 4'h0;
assign strg_ub_agg_read_addr_gen_0_strides_3 = 8'h0;
assign strg_ub_agg_read_addr_gen_0_strides_4 = 8'h0;
assign strg_ub_agg_read_addr_gen_0_strides_5 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_strides_0 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_strides_1 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_strides_2 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_strides_3 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_strides_4 = 8'h0;
assign strg_ub_agg_read_addr_gen_1_strides_5 = 8'h0;
assign strg_ub_tb_write_addr_gen_1_starting_addr_0 = 6'h0;
assign strg_ub_tb_write_addr_gen_1_starting_addr_1 = 6'h0;
assign strg_ub_tb_write_addr_gen_1_starting_addr_2 = 6'h0;
assign strg_ub_tb_write_addr_gen_1_starting_addr_3 = 6'h0;
assign strg_ub_tb_write_addr_gen_1_starting_addr_4 = 6'h0;
assign strg_ub_tb_write_addr_gen_1_starting_addr_5 = 6'h0;
assign strg_ub_output_addr_gen_starting_addr_0 = 16'h0;
assign strg_ub_output_addr_gen_starting_addr_1 = 16'h0;
assign strg_ub_output_addr_gen_starting_addr_2 = 16'h0;
assign strg_ub_output_addr_gen_starting_addr_3 = 16'h0;
assign strg_ub_output_addr_gen_starting_addr_4 = 16'h0;
assign strg_ub_output_addr_gen_starting_addr_5 = 16'h0;
assign strg_ub_tb_write_addr_gen_1_strides_4 = 6'h0;
assign strg_ub_tb_write_addr_gen_1_strides_5 = 6'h0;
assign strg_ub_tb_write_addr_gen_0_starting_addr_0 = 6'h0;
assign strg_ub_tb_write_addr_gen_0_starting_addr_1 = 6'h0;
assign strg_ub_tb_write_addr_gen_0_starting_addr_2 = 6'h0;
assign strg_ub_tb_write_addr_gen_0_starting_addr_3 = 6'h0;
assign strg_ub_tb_write_addr_gen_0_starting_addr_4 = 6'h0;
assign strg_ub_tb_write_addr_gen_0_starting_addr_5 = 6'h0;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality_0 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality_1 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality_2 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality_3 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality_4 = 3'h0;
assign strg_ub_loops_in2buf_autovec_read_0_dimensionality_5 = 3'h0;
assign strg_ub_agg_write_addr_gen_1_strides_0 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_strides_1 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_strides_2 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_strides_3 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_strides_4 = 4'h0;
assign strg_ub_agg_write_addr_gen_1_strides_5 = 4'h0;
assign strg_ub_output_addr_gen_strides_4 = 16'h0;
assign strg_ub_output_addr_gen_strides_5 = 16'h0;
assign strg_ub_loops_in2buf_autovec_read_1_ranges_0 = 8'h0;
assign strg_ub_loops_in2buf_autovec_read_1_ranges_1 = 8'h0;
assign strg_ub_loops_in2buf_autovec_read_1_ranges_2 = 8'h0;
assign strg_ub_loops_in2buf_autovec_read_1_ranges_3 = 8'h0;
assign strg_ub_loops_in2buf_autovec_read_1_ranges_4 = 8'h0;
assign strg_ub_loops_in2buf_autovec_read_1_ranges_5 = 8'h0;
assign strg_ub_agg_write_addr_gen_0_starting_addr_0 = 4'h0;
assign strg_ub_agg_write_addr_gen_0_starting_addr_1 = 4'h0;
assign strg_ub_agg_write_addr_gen_0_starting_addr_2 = 4'h0;
assign strg_ub_agg_write_addr_gen_0_starting_addr_3 = 4'h0;
assign strg_ub_agg_write_addr_gen_0_starting_addr_4 = 4'h0;
assign strg_ub_agg_write_addr_gen_0_starting_addr_5 = 4'h0;
assign strg_ub_loops_in2buf_1_ranges_0 = 4'h0;
assign strg_ub_loops_in2buf_1_ranges_1 = 4'h0;
assign strg_ub_loops_in2buf_1_ranges_2 = 4'h0;
assign strg_ub_loops_in2buf_1_ranges_3 = 4'h0;
assign strg_ub_loops_in2buf_1_ranges_4 = 4'h0;
assign strg_ub_loops_in2buf_1_ranges_5 = 4'h0;
assign strg_ub_input_addr_gen_strides_3 = 16'h0;
assign strg_ub_input_addr_gen_strides_4 = 16'h0;
assign strg_ub_input_addr_gen_strides_5 = 16'h0;
assign strg_ub_out_port_sel_addr_starting_addr_0 = 1'h0;
assign strg_ub_out_port_sel_addr_starting_addr_1 = 1'h0;
assign strg_ub_out_port_sel_addr_starting_addr_2 = 1'h0;
assign strg_ub_out_port_sel_addr_starting_addr_3 = 1'h0;
assign strg_ub_out_port_sel_addr_starting_addr_4 = 1'h0;
assign strg_ub_out_port_sel_addr_starting_addr_5 = 1'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr_0 = 16'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr_1 = 16'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr_2 = 16'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr_3 = 16'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr_4 = 16'h0;
assign strg_ub_tb_read_sched_gen_1_sched_addr_gen_starting_addr_5 = 16'h0;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality_0 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality_1 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality_2 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality_3 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality_4 = 2'h0;
assign strg_ub_loops_buf2out_autovec_write_1_dimensionality_5 = 2'h0;
assign strg_ub_tb_read_addr_gen_1_starting_addr_0 = 6'h0;
assign strg_ub_tb_read_addr_gen_1_starting_addr_1 = 6'h0;
assign strg_ub_tb_read_addr_gen_1_starting_addr_2 = 6'h0;
assign strg_ub_tb_read_addr_gen_1_starting_addr_3 = 6'h0;
assign strg_ub_tb_read_addr_gen_1_starting_addr_4 = 6'h0;
assign strg_ub_tb_read_addr_gen_1_starting_addr_5 = 6'h0;
assign strg_ub_loops_buf2out_read_1_dimensionality_0 = 2'h0;
assign strg_ub_loops_buf2out_read_1_dimensionality_1 = 2'h0;
assign strg_ub_loops_buf2out_read_1_dimensionality_2 = 2'h0;
assign strg_ub_loops_buf2out_read_1_dimensionality_3 = 2'h0;
assign strg_ub_loops_buf2out_read_1_dimensionality_4 = 2'h0;
assign strg_ub_loops_buf2out_read_1_dimensionality_5 = 2'h0;
assign strg_ub_tb_write_addr_gen_0_strides_4 = 6'h0;
assign strg_ub_tb_write_addr_gen_0_strides_5 = 6'h0;

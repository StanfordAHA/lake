`timescale 1ns/1ns
`ifndef TX_NUM_GLB
`define TX_NUM_GLB 1
`endif

module vector_reducer_tb;

    reg clk;
    reg clk_en;
    reg rst_n;
    reg stall;
    reg flush;
    reg tile_en;
    reg vector_reduce_mode;
    reg joiner_op; 
    wire [63:0] cycle_count ;

    // wire for dut input & output
    wire [16:0] crddrp_crd_in;
    wire crddrp_crd_in_valid;
    wire crddrp_crd_in_ready;

    wire [16:0] mult_val_in;
    wire mult_val_in_valid;
    wire mult_val_in_ready;

    wire [16:0] read_scanner_ext_us_pos_in;
    wire read_scanner_ext_us_pos_in_valid;
    wire read_scanner_ext_us_pos_in_ready;

    wire [16:0] final_column_coords_out;
    wire final_column_coords_out_valid;
    wire final_column_coords_out_ready;

    wire [16:0] final_vals_out;
    wire final_vals_out_valid;
    wire final_vals_out_ready;

    wire [16:0] coord_out;
    wire coord_out_valid;
    wire coord_out_ready;

    wire [16:0] union_val_out_0;
    wire union_val_out_0_valid;

    wire [16:0] union_val_out_1;
    wire union_val_out_1_valid;

    wire [16:0] loop_val_out;
    wire loop_val_out_ready;

    wire [16:0] loop_column_coords_out;
    wire loop_column_coords_out_ready;
    wire loop_column_coords_out_valid;

    wire [16:0] loop_column_coords_in;
    wire loop_column_coords_in_ready;
    wire loop_column_coords_in_valid;

    wire [16:0] loop_vals_in;
    wire loop_vals_in_ready;
    wire loop_vals_in_valid;

    // wire for mem
    wire [63:0] memory_0_data_in_p0;
    wire [63:0] memory_0_data_out_p0;
    wire [8:0] memory_addr_to_mem_p0;
    wire memory_0_read_enable_p0;
    wire memory_0_write_enable_p0;

    wire [63:0] memory_1_data_in_p1;
    wire [63:0] memory_1_data_out_p1;
    wire [8:0] memory_addr_to_mem_p1;
    wire memory_1_read_enable_p1;
    wire memory_1_write_enable_p1;

    // dummy connection
    wire [16:0] ws_addr;
    wire ws_addr_valid;
    wire ws_addr_ready;

    wire [16:0] ws_blk;
    wire ws_blk_valid;
    wire ws_blk_ready;

    wire [16:0] rs_blk;
    wire rs_blk_valid;
    wire rs_blk_ready;

    assign {ws_addr, ws_addr_valid, ws_blk, ws_blk_valid} = 35'b0;
    assign {rs_blk, rs_blk_valid} = 17'b0;

    logic [1:0] [31:0] config_out;

    wire [4:0] done;
    parameter NUM_CYCLES = 40000;

    integer clk_count;
    integer start_write;
    integer write_eos;
    integer write_count;
    logic start_read;
    logic read_input_in;
    integer read_count;
    integer wait_gap = 0; // should pass with arb gap
    integer DONE_TOKEN = 17'h10100;

    intersect_unit #(    
    ) dut (
        .clk(clk),
        .clk_en(clk_en),
        .coord_in_0(crddrp_crd_in),
        .coord_in_0_valid(crddrp_crd_in_valid),
        .coord_in_0_ready(crddrp_crd_in_ready),
        .coord_in_1(loop_column_coords_in),
        .coord_in_1_valid(loop_column_coords_in_valid),
        .coord_in_1_ready(loop_column_coords_in_ready),
        .pos_in_0(mult_val_in),
        .pos_in_0_valid(mult_val_in_valid),
        .pos_in_0_ready(mult_val_in_ready),
        .pos_in_1(loop_vals_in),
        .pos_in_1_valid(loop_vals_in_valid),
        .pos_in_1_ready(loop_vals_in_ready),
        .joiner_op(joiner_op),
        .tile_en(tile_en),
        .coord_out(loop_column_coords_out),
        .coord_out_valid(loop_column_coords_out_valid),
        .coord_out_ready(loop_column_coords_out_ready),
        .pos_out_0(union_val_out_0),
        .pos_out_0_valid(union_val_out_0_valid),
        .pos_out_0_ready(loop_val_out_ready),
        .pos_out_1(union_val_out_1),
        .pos_out_1_valid(union_val_out_1_valid),
        .pos_out_1_ready(loop_val_out_ready),
        .rst_n(rst_n),
        .flush(flush),
        .tile_en(tile_en),
        .vector_reduce_mode(vector_reduce_mode)
    );

    fiber_access_16 fiber_access_coords 
    (
    .buffet_buffet_capacity_log({4'b1000, 4'b1000}),
    .data_from_mem(memory_0_data_out_p0),
    .buffet_tile_en(tile_en),
    .clk(clk),
    .clk_en(clk_en),
    .flush(flush),
    .read_scanner_block_mode(1'b0),
    .read_scanner_block_rd_out_ready(rs_blk_ready),
    .read_scanner_coord_out_ready(loop_column_coords_in_ready),
    .read_scanner_dense(1'b0),
    .read_scanner_dim_size(16'b0),
    .read_scanner_do_repeat(1'b0),
    .read_scanner_inner_dim_offset(16'b0),
    .read_scanner_lookup(1'b0),
    .read_scanner_pos_out_ready(final_column_coords_out_ready),
    .read_scanner_repeat_factor(16'b0),
    .read_scanner_repeat_outer_inner_n(1'b0),
    .read_scanner_root(1'b0),
    // .read_scanner_spacc_mode(1'b0),
    // .read_scanner_stop_lvl(16'b0),
    .read_scanner_tile_en(tile_en),
    .read_scanner_us_pos_in(read_scanner_ext_us_pos_in),
    // .read_scanner_us_pos_in_valid(pos_in_0_valid & start_read == 1),
    .read_scanner_us_pos_in_valid(read_scanner_ext_us_pos_in_valid),
    .rst_n(rst_n),
    .tile_en(tile_en),
    .write_scanner_addr_in(ws_addr),
    .write_scanner_addr_in_valid(ws_addr_valid),
    .write_scanner_block_mode(1'b0),
    .write_scanner_block_wr_in(ws_blk),
    .write_scanner_block_wr_in_valid(ws_blk_valid),
    .write_scanner_compressed(1'b1),
    .write_scanner_data_in(loop_column_coords_out),
    .write_scanner_data_in_valid(loop_column_coords_out_valid),
    .write_scanner_init_blank(1'b0),
    .write_scanner_lowest_level(1'b0),
    // .write_scanner_spacc_mode(1'b0),
    // .write_scanner_stop_lvl(16'b0),
    .write_scanner_tile_en(tile_en),
    .addr_to_mem(memory_addr_to_mem_p0),
    .data_to_mem(memory_0_data_in_p0),
    .read_scanner_block_rd_out(rs_blk),
    .read_scanner_block_rd_out_valid(rs_blk_valid),
    .read_scanner_coord_out(loop_column_coords_in),
    .read_scanner_coord_out_valid(loop_column_coords_in_valid),
    .read_scanner_pos_out(final_column_coords_out),
    .read_scanner_pos_out_valid(final_column_coords_out_valid),
    .read_scanner_us_pos_in_ready(read_scanner_ext_us_pos_in_ready),
    .ren_to_mem(memory_0_read_enable_p0),
    .wen_to_mem(memory_0_write_enable_p0),
    .write_scanner_addr_in_ready(ws_addr_ready),
    .write_scanner_block_wr_in_ready(ws_blk_ready),
    .write_scanner_data_in_ready(loop_column_coords_out_ready),
    .vector_reduce_mode(vector_reduce_mode)
    );


    fiber_access_16 fiber_access_vals 
    (
    .buffet_buffet_capacity_log({4'b1000, 4'b1000}),
    .data_from_mem(memory_1_data_out_p1),
    .buffet_tile_en(tile_en),
    .clk(clk),
    .clk_en(clk_en),
    .flush(flush),
    .read_scanner_block_mode(1'b0),
    .read_scanner_block_rd_out_ready(rs_blk_ready),
    .read_scanner_coord_out_ready(loop_vals_in_ready),
    .read_scanner_dense(1'b0),
    .read_scanner_dim_size(16'b0),
    .read_scanner_do_repeat(1'b0),
    .read_scanner_inner_dim_offset(16'b0),
    .read_scanner_lookup(1'b0),
    .read_scanner_pos_out_ready(final_vals_out_ready),
    .read_scanner_repeat_factor(16'b0),
    .read_scanner_repeat_outer_inner_n(1'b0),
    .read_scanner_root(1'b0),
    // .read_scanner_spacc_mode(1'b0),
    // .read_scanner_stop_lvl(16'b0),
    .read_scanner_tile_en(tile_en),
    .read_scanner_us_pos_in(read_scanner_ext_us_pos_in),
    // .read_scanner_us_pos_in_valid(pos_in_0_valid & start_read == 1),
    .read_scanner_us_pos_in_valid(read_scanner_ext_us_pos_in_valid),
    .rst_n(rst_n),
    .tile_en(tile_en),
    .write_scanner_addr_in(ws_addr),
    .write_scanner_addr_in_valid(ws_addr_valid),
    .write_scanner_block_mode(1'b0),
    .write_scanner_block_wr_in(ws_blk),
    .write_scanner_block_wr_in_valid(ws_blk_valid),
    .write_scanner_compressed(1'b1),
    .write_scanner_data_in(loop_val_out),
    .write_scanner_data_in_valid(union_val_out_0_valid & union_val_out_1_valid), // PAY ATTENTION TO THIS
    .write_scanner_init_blank(1'b0),
    .write_scanner_lowest_level(1'b0),
    // .write_scanner_spacc_mode(1'b0),
    // .write_scanner_stop_lvl(16'b0),
    .write_scanner_tile_en(tile_en),
    .addr_to_mem(memory_addr_to_mem_p1),
    .data_to_mem(memory_1_data_in_p1),
    .read_scanner_block_rd_out(rs_blk),
    .read_scanner_block_rd_out_valid(rs_blk_valid),
    .read_scanner_coord_out(loop_vals_in),
    .read_scanner_coord_out_valid(loop_vals_in_valid),
    .read_scanner_pos_out(final_vals_out),
    .read_scanner_pos_out_valid(final_vals_out_valid),
    .read_scanner_us_pos_in_ready(read_scanner_ext_us_pos_in_ready),
    .ren_to_mem(memory_1_read_enable_p1),
    .wen_to_mem(memory_1_write_enable_p1),
    .write_scanner_addr_in_ready(ws_addr_ready),
    .write_scanner_block_wr_in_ready(ws_blk_ready),
    .write_scanner_data_in_ready(loop_val_out_ready),
    .vector_reduce_mode(vector_reduce_mode)
    );

    behavioral_pe_add behavioral_pe_add
    (
        .a_in(union_val_out_0),
        .b_in(union_val_out_1),
        .out(loop_val_out)
    );

    glb_write #(
        .FILE_NAME("crddrp_crd_in.txt"),
        .TX_NUM(`TX_NUM_GLB),
        .RAN_SHITF(0)
    ) crddrp_crd_in_inst (
        .clk(clk),
        .rst_n(rst_n),
        .data(crddrp_crd_in),
        // .ready(pos_in_0_ready & start_read == 1),
        .ready(crddrp_crd_in_ready),
        .valid(crddrp_crd_in_valid),
        .done(done[0]),
        .flush(flush)
    );

    glb_write #(
        .FILE_NAME("mult_val_in.txt"),
        .TX_NUM(`TX_NUM_GLB),
        .RAN_SHITF(0)
    ) mult_val_in_inst (
        .clk(clk),
        .rst_n(rst_n),
        .data(mult_val_in),
        .ready(mult_val_in_ready),
        .valid(mult_val_in_valid),
        .done(done[1]),
        .flush(flush)
    );

    // DUMMY 
    glb_write #(
        .FILE_NAME("ext_us_pos_in.txt"),
        .TX_NUM(`TX_NUM_GLB),
        .RAN_SHITF(0)
    ) fiber_access_ext_us_pos_in_inst (
        .clk(clk),
        .rst_n(rst_n),
        .data(read_scanner_ext_us_pos_in),
        // .ready(pos_in_0_ready & start_read == 1),
        .ready(read_scanner_ext_us_pos_in_ready),
        .valid(read_scanner_ext_us_pos_in_valid),
        .done(done[2]),
        .flush(flush)
    );

    glb_read #(
        .FILE_NAME("column_coords_out.txt"),
        .TX_NUM(`TX_NUM_GLB),
        .RAN_SHITF(0)
    ) final_column_coords_out_inst (
        .clk(clk),
        .rst_n(rst_n),
        .data(final_column_coords_out),
        .ready(final_column_coords_out_ready),
        .valid(final_column_coords_out_valid),
        .done(done[3]),
        .flush(flush)
    );

    glb_read #(
        .FILE_NAME("vals_out.txt"),
        .TX_NUM(`TX_NUM_GLB),
        .RAN_SHITF(0)
    ) final_vals_out_inst (
        .clk(clk),
        .rst_n(rst_n),
        .data(final_vals_out),
        .ready(final_vals_out_ready),
        .valid(final_vals_out_valid),
        .done(done[4]),
        .flush(flush)
    );

    sram_sp memory_0 (
        .clk(clk),
        .clk_en(clk_en),
        .data_in_p0(memory_0_data_in_p0),
        .flush(flush),
        .read_addr_p0(memory_addr_to_mem_p0),
        .read_enable_p0(memory_0_read_enable_p0),
        .write_addr_p0(memory_addr_to_mem_p0),
        .write_enable_p0(memory_0_write_enable_p0),
        .data_out_p0(memory_0_data_out_p0)
    );


    sram_sp memory_1 (
        .clk(clk),
        .clk_en(clk_en),
        .data_in_p0(memory_1_data_in_p1),
        .flush(flush),
        .read_addr_p0(memory_addr_to_mem_p1),
        .read_enable_p0(memory_1_read_enable_p1),
        .write_addr_p0(memory_addr_to_mem_p1),
        .write_enable_p0(memory_1_write_enable_p1),
        .data_out_p0(memory_1_data_out_p1)
    );

    // simulated clk signal, 10ns period
    initial begin
        clk_count = 0;
        start_write = 0;
        write_eos = 0;
        write_count = 0;
        start_read = 0;
        read_input_in = 0;
        read_count = 0;

        clk = 0;
        clk_en = 1;
        rst_n = 0;
        tile_en = 1;
        joiner_op = 1;
        vector_reduce_mode = 1;
        flush = 0;

        #5 clk = 1;
        flush = 1;
        rst_n = 1;
        #5 clk = 0;
        flush = 0;

        for(integer i = 0; i < NUM_CYCLES * 2; i = i + 1) begin
            #5 clk = ~clk;

        end
        //$display("write cycle count: %0d", write_count);
        //$display("read cycle count: %0d", read_count);
        $finish;
    
    end

endmodule
